LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY mux_3bits IS
    PORT (
        IN1, IN2, IN3, IN4, IN5 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        SEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
        SELECTED : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE arch_mux_3bits OF mux_3bits IS
BEGIN
    SELECTED <= IN1 WHEN sel = "000" ELSE
        IN2 WHEN SEL = "001" ELSE
        IN3 WHEN SEL = "010" ELSE
        IN4 WHEN SEL = "011" ELSE
        IN5 WHEN SEL = "100";
END ARCHITECTURE;
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE std.STANDARD.NATURAL;
USE ieee.numeric_std.ALL;
--Entity B
ENTITY alu IS
    PORT (
        src1, src2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        ALU_signal : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
        result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
        flags : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE arch_alu OF alu IS
    SIGNAL one : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL zero : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL temp : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
    zero <= (OTHERS => '0');
    one <= (0 => '1', OTHERS => '0');
    temp <= (to_integer(unsigned(src2)) => '1', OTHERS => '0');

    result <= NOT src2 WHEN ALU_signal = "0001" ELSE
        zero - src2 WHEN ALU_signal = "0010" ELSE
        src2 + one WHEN ALU_signal = "0011" ELSE
        src2 - one WHEN ALU_signal = "0100" ELSE
        src1 + src2 WHEN ALU_signal = "0110" ELSE
        src1 - src2 WHEN ALU_signal = "0111" ELSE
        src1 AND src2 WHEN ALU_signal = "1000" ELSE
        src1 OR src2 WHEN ALU_signal = "1001" ELSE
        src1 XOR src2 WHEN ALU_signal = "1010" ELSE
        src1 OR temp WHEN ALU_signal = "1011" ELSE
        src2(0) & src2(31 DOWNTO 1) WHEN ALU_signal = "1101" ELSE
        src2(30 DOWNTO 0) & src2(31) WHEN ALU_signal = "1100";

END ARCHITECTURE;
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY mux_3bits IS
    PORT (
        IN1, IN2, IN3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        SEL : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
        SELECTED : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE arch_mux_3bits OF mux_3bits IS
BEGIN
    SELECTED <= IN1 WHEN sel = "00" ELSE
        IN2 WHEN SEL = "01" ELSE
        IN3 WHEN SEL = "10";
END ARCHITECTURE;